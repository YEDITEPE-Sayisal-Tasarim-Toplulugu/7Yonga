


`ifndef __SOC_CINFIGURATION_SVH__
`define __SOC_CINFIGURATION_SVH__

package soc_config_pkg;

// Parametrik sabitler
parameter int USE_SOFT_MEMORY_MODULES = 1;
parameter int USE_SOFT_ROM_MODULES = 1;

endpackage

`endif // __SOC_CINFIGURATION_SVH__