`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 16.05.2025 21:10:25
// Design Name: 
// Module Name: soc_peripherals_top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module soc_peripherals_top
    #(
    )
    (
        input logic clk_i, reset_i,
        
        AXI_BUS.Slave              AXI4_slave
    );
    
    
    
endmodule













