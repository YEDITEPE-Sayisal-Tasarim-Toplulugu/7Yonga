// Copyright 2025 Yeditepe Üniversitesi Sayısal Tasarım Topluluğu.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.

////////////////////////////////////////////////////////////////////////////////
// Engineer:       M. Furkan UZUN - @mfu                                      //
//                                                                            //
//                                                                            //
// Design Name:    CV32E40P Instruction and Data Memory Interfaces            //
// Project Name:   7Yonga                                                     //
// Language:       SystemVerilog                                              //
//                                                                            //
// Description:    CV32E40P Instruction and Data Memory Interfaces tanımları  //
//                                                                            //
////////////////////////////////////////////////////////////////////////////////

`ifndef __SOC_INTERFACE_LIST_SVH__
`define __SOC_INTERFACE_LIST_SVH__

interface CV32E_INST_INF();
    logic [31:0] instr_addr;
    logic instr_req;
    logic instr_gnt;
    logic instr_rvalid;
    logic [31:0] instr_rdata;
    
    modport MASTER
    (
        output instr_addr,
        output instr_req,
        input instr_gnt,
        input instr_rvalid,
        input instr_rdata
    );
    
    modport SLAVE
    (
        input instr_addr,
        input instr_req,
        output instr_gnt,
        output instr_rvalid,
        output instr_rdata
    );
    
endinterface


interface CV32E_DATA_INF();
    logic [31:0] data_addr;
    logic data_req;
    logic data_gnt;
    logic data_we;
    logic [3:0] data_be;
    logic [31:0] data_wdata;
    logic data_rvalid;
    logic [31:0] data_rdata;
    
    modport MASTER
    (
        output data_addr,
        output data_req,
        input data_gnt,
        output data_we,
        output data_be,
        output data_wdata,
        input data_rvalid,
        input data_rdata
    );
    
    modport SLAVE
    (
        input data_addr,
        input data_req,
        output data_gnt,
        input data_we,
        input data_be,
        input data_wdata,
        output data_rvalid,
        output data_rdata
    );
    
endinterface

`endif //__SOC_INTERFACE_LIST_SVH__










